//switched to wordirbranch
module top.v (
	input  clk_i,
	input  rst_i,
	input  a_i,
	output z_o
);

assign z_o = a_i;
endmodule
